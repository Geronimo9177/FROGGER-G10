/*######################################################################
//#	G0B1T: HDL EXAMPLES. 2018.
//######################################################################
//# Copyright (C) 2018. F.E.Segura-Quijano (FES) fsegura@uniandes.edu.co
//# 
//# This program is free software: you can redistribute it and/or modify
//# it under the terms of the GNU General Public License as published by
//# the Free Software Foundation, version 3 of the License.
//#
//# This program is distributed in the hope that it will be useful,
//# but WITHOUT ANY WARRANTY; without even the implied warranty of
//# MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//# GNU General Public License for more details.
//#
//# You should have received a copy of the GNU General Public License
//# along with this program.  If not, see <http://www.gnu.org/licenses/>
//####################################################################*/
//=======================================================
//  MODULE Definition
//=======================================================
module SC_LEVELCOUNTER (
	//////////// OUTPUTS //////////
	SC_LEVEL_COUNTER_data_OutBUS,
	//////////// INPUTS //////////
	SC_LEVEL_COUNTER_CLOCK_50,
	SC_LEVEL_COUNTER_RESET_InHigh,
	SC_LEVEL_COUNTER_CUENTA_InLow
);
//=======================================================
//  PARAMETER declarations
//=======================================================
parameter DATAWIDTH_3 = 3;
//=======================================================
//  PORT declarations
//=======================================================
output	[DATAWIDTH_3-1:0]	SC_LEVEL_COUNTER_data_OutBUS;
input		SC_LEVEL_COUNTER_CLOCK_50;
input		SC_LEVEL_COUNTER_RESET_InHigh;
input		[DATAWIDTH_3-1:0] SC_LEVEL_COUNTER_CUENTA_InLow;
//=======================================================
//  REG/WIRE declarations
//=======================================================
reg [DATAWIDTH_3-1:0] LEVELCOUNTER_Register;
reg [DATAWIDTH_3-1:0] LEVELCOUNTER_Signal;
//=======================================================
//  Structural coding
//=======================================================
//INPUT LOGIC: COMBINATIONAL
always @(*)
begin
	if (SC_LEVEL_COUNTER_CUENTA_InLow == 3'b000)
		LEVELCOUNTER_Signal = LEVELCOUNTER_Register + 1'b1;
	else if (SC_LEVEL_COUNTER_CUENTA_InLow == 3'b111)
		LEVELCOUNTER_Signal = LEVELCOUNTER_Register;
	else
		LEVELCOUNTER_Signal = SC_LEVEL_COUNTER_CUENTA_InLow;
	end	
//STATE REGISTER: SEQUENTIAL
always @(posedge SC_LEVEL_COUNTER_CLOCK_50, posedge SC_LEVEL_COUNTER_RESET_InHigh)
begin
	if (SC_LEVEL_COUNTER_RESET_InHigh == 1'b1)
		LEVELCOUNTER_Register <= 3'b001;
	else
		LEVELCOUNTER_Register <= LEVELCOUNTER_Signal;
end
//=======================================================
//  Outputs
//=======================================================
//OUTPUT LOGIC: COMBINATIONAL
assign SC_LEVEL_COUNTER_data_OutBUS = LEVELCOUNTER_Register;

endmodule
