/*######################################################################
//#	G0B1T: HDL EXAMPLES. 2018.
//######################################################################
//# Copyright (C) 2018. F.E.Segura-Quijano (FES) fsegura@uniandes.edu.co
//# 
//# This program is free software: you can redistribute it and/or modify
//# it under the terms of the GNU General Public License as published by
//# the Free Software Foundation, version 3 of the License.
//#
//# This program is distributed in the hope that it will be useful,
//# but WITHOUT ANY WARRANTY; without even the implied warranty of
//# MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//# GNU General Public License for more details.
//#
//# You should have received a copy of the GNU General Public License
//# along with this program.  If not, see <http://www.gnu.org/licenses/>
//####################################################################*/
//=======================================================
//  MODULE Definition
//=======================================================
module SC_LIFECOUNTER (
	//////////// OUTPUTS //////////
	SC_LIFE_COUNTER_data_OutBUS,
	//////////// INPUTS //////////
	SC_LIFE_COUNTER_CLOCK_50,
	SC_LIFE_COUNTER_RESET_InHigh,
	SC_LIFE_COUNTER_CUENTA_InLow
);
//=======================================================
//  PARAMETER declarations
//=======================================================
parameter DATAWIDTH_2 = 2;
//=======================================================
//  PORT declarations
//=======================================================
output	[DATAWIDTH_2-1:0]	SC_LIFE_COUNTER_data_OutBUS;
input		SC_LIFE_COUNTER_CLOCK_50;
input		SC_LIFE_COUNTER_RESET_InHigh;
input		SC_LIFE_COUNTER_CUENTA_InLow;
//=======================================================
//  REG/WIRE declarations
//=======================================================
reg [DATAWIDTH_2-1:0] LIFECOUNTER_Register;
reg [DATAWIDTH_2-1:0] LIFECOUNTER_Signal;
//=======================================================
//  Structural coding
//=======================================================
//INPUT LOGIC: COMBINATIONAL
always @(*)
begin
	if (SC_LIFE_COUNTER_CUENTA_InLow == 1'b0)
		LIFECOUNTER_Signal = LIFECOUNTER_Register - 1'b1;
	else
		LIFECOUNTER_Signal = LIFECOUNTER_Register;
	end	
//STATE REGISTER: SEQUENTIAL
always @(posedge SC_LIFE_COUNTER_CLOCK_50, posedge SC_LIFE_COUNTER_RESET_InHigh)
begin
	if (SC_LIFE_COUNTER_RESET_InHigh == 1'b1)
		LIFECOUNTER_Register <= 2'b11;
	else
		LIFECOUNTER_Register <= LIFECOUNTER_Signal;
end
//=======================================================
//  Outputs
//=======================================================
//OUTPUT LOGIC: COMBINATIONAL
assign SC_LIFE_COUNTER_data_OutBUS = LIFECOUNTER_Register;

endmodule
