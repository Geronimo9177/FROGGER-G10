/*######################################################################
//#	G0B1T: HDL EXAMPLES. 2018.
//######################################################################
//# Copyright (C) 2018. F.E.Segura-Quijano (FES) fsegura@uniandes.edu.co
//# 
//# This program is free software: you can redistribute it and/or modify
//# it under the terms of the GNU General Public License as published by
//# the Free Software Foundation, version 3 of the License.
//#
//# This program is distributed in the hope that it will be useful,
//# but WITHOUT ANY WARRANTY; without even the implied warranty of
//# MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//# GNU General Public License for more details.
//#
//# You should have received a copy of the GNU General Public License
//# along with this program.  If not, see <http://www.gnu.org/licenses/>
//####################################################################*/
//=======================================================
//  MODULE Definition
//=======================================================
module CC_COMPARATORCRASH (
//////////// OUTPUTS //////////
	CC_COMPARADORCRASH_Out_Bus,
	CC_COMPARATORLOCATION_Out,
//////////// INPUTS //////////
	CC_COMPARADORCRASH_ALBERT_FROG_ROW_2_In_Bus,
	CC_COMPARADORCRASH_ALBERT_FROG_ROW_3_In_Bus,
	CC_COMPARADORCRASH_ALBERT_FROG_ROW_4_In_Bus,
	CC_COMPARADORCRASH_ALBERT_FROG_ROW_5_In_Bus,
	CC_COMPARADORCRASH_ALBERT_FROG_ROW_6_In_Bus,
	CC_COMPARADORCRASH_ALBERT_FROG_ROW_7_In_Bus,
	CC_COMPARADORCRASH_ALBERT_FROG_ROW_8_In_Bus,
	CC_COMPARADORCRASH_ALBERT_FROG_ROW_9_In_Bus,
	CC_COMPARADORCRASH_ALBERT_FROG_ROW_10_In_Bus,
	CC_COMPARADORCRASH_ALBERT_FROG_ROW_11_In_Bus,
	CC_COMPARADORCRASH_ALBERT_FROG_ROW_12_In_Bus,
	CC_COMPARADORCRASH_ALBERT_FROG_ROW_13_In_Bus,
	CC_COMPARADORCRASH_ALBERT_FROG_ROW_14_In_Bus,

	CC_COMPARADORCRASH_BACKGROUND_ROW_2_IN_BUS,
	CC_COMPARADORCRASH_BACKGROUND_ROW_3_IN_BUS,
	CC_COMPARADORCRASH_BACKGROUND_ROW_4_IN_BUS,
	CC_COMPARADORCRASH_BACKGROUND_ROW_5_IN_BUS,
	CC_COMPARADORCRASH_BACKGROUND_ROW_6_IN_BUS,
	CC_COMPARADORCRASH_BACKGROUND_ROW_9_IN_BUS,
	CC_COMPARADORCRASH_BACKGROUND_ROW_10_IN_BUS,
	CC_COMPARADORCRASH_BACKGROUND_ROW_11_IN_BUS,
	CC_COMPARADORCRASH_BACKGROUND_ROW_12_IN_BUS,
	CC_COMPARADORCRASH_BACKGROUND_ROW_13_IN_BUS,
	CC_COMPARADORCRASH_END_GOAL_ROW_14_IN_BUS,
	
	CC_COMPARADORCRASH_IMAGE_INBUS
);
//=======================================================
//  PARAMETER declarations
//=======================================================
parameter DATAWIDTH_BUS = 8;
parameter DATAWIDTH_OUT_BUS = 2;
//=======================================================
//  PORT declarations
//=======================================================
output	reg [DATAWIDTH_OUT_BUS-1:0] CC_COMPARADORCRASH_Out_Bus;
output	reg CC_COMPARATORLOCATION_Out;
input 	[DATAWIDTH_BUS-1:0] CC_COMPARADORCRASH_ALBERT_FROG_ROW_2_In_Bus;
input 	[DATAWIDTH_BUS-1:0] CC_COMPARADORCRASH_ALBERT_FROG_ROW_3_In_Bus;
input 	[DATAWIDTH_BUS-1:0] CC_COMPARADORCRASH_ALBERT_FROG_ROW_4_In_Bus;
input 	[DATAWIDTH_BUS-1:0] CC_COMPARADORCRASH_ALBERT_FROG_ROW_5_In_Bus;
input 	[DATAWIDTH_BUS-1:0] CC_COMPARADORCRASH_ALBERT_FROG_ROW_6_In_Bus;
input 	[DATAWIDTH_BUS-1:0] CC_COMPARADORCRASH_ALBERT_FROG_ROW_7_In_Bus;
input 	[DATAWIDTH_BUS-1:0] CC_COMPARADORCRASH_ALBERT_FROG_ROW_8_In_Bus;
input 	[DATAWIDTH_BUS-1:0] CC_COMPARADORCRASH_ALBERT_FROG_ROW_9_In_Bus;
input 	[DATAWIDTH_BUS-1:0] CC_COMPARADORCRASH_ALBERT_FROG_ROW_10_In_Bus;
input 	[DATAWIDTH_BUS-1:0] CC_COMPARADORCRASH_ALBERT_FROG_ROW_11_In_Bus;
input 	[DATAWIDTH_BUS-1:0] CC_COMPARADORCRASH_ALBERT_FROG_ROW_12_In_Bus;
input 	[DATAWIDTH_BUS-1:0] CC_COMPARADORCRASH_ALBERT_FROG_ROW_13_In_Bus;
input 	[DATAWIDTH_BUS-1:0] CC_COMPARADORCRASH_ALBERT_FROG_ROW_14_In_Bus;
input 	[DATAWIDTH_BUS-1:0] CC_COMPARADORCRASH_BACKGROUND_ROW_2_IN_BUS;
input 	[DATAWIDTH_BUS-1:0] CC_COMPARADORCRASH_BACKGROUND_ROW_3_IN_BUS;
input 	[DATAWIDTH_BUS-1:0] CC_COMPARADORCRASH_BACKGROUND_ROW_4_IN_BUS;
input 	[DATAWIDTH_BUS-1:0] CC_COMPARADORCRASH_BACKGROUND_ROW_5_IN_BUS;
input 	[DATAWIDTH_BUS-1:0] CC_COMPARADORCRASH_BACKGROUND_ROW_6_IN_BUS;
input 	[DATAWIDTH_BUS-1:0] CC_COMPARADORCRASH_BACKGROUND_ROW_9_IN_BUS;
input 	[DATAWIDTH_BUS-1:0] CC_COMPARADORCRASH_BACKGROUND_ROW_10_IN_BUS;
input 	[DATAWIDTH_BUS-1:0] CC_COMPARADORCRASH_BACKGROUND_ROW_11_IN_BUS;
input 	[DATAWIDTH_BUS-1:0] CC_COMPARADORCRASH_BACKGROUND_ROW_12_IN_BUS;
input 	[DATAWIDTH_BUS-1:0] CC_COMPARADORCRASH_BACKGROUND_ROW_13_IN_BUS;
input 	[DATAWIDTH_BUS-1:0] CC_COMPARADORCRASH_END_GOAL_ROW_14_IN_BUS;
input    [1:0] CC_COMPARADORCRASH_IMAGE_INBUS;

//=======================================================
//  REG/WIRE declarations
//=======================================================
//=======================================================
//  Structural coding
//=======================================================
always @(*)
begin
	if (CC_COMPARADORCRASH_IMAGE_INBUS == 2'b10)
		CC_COMPARADORCRASH_Out_Bus = 2'b00;
	else if ((CC_COMPARADORCRASH_ALBERT_FROG_ROW_2_In_Bus != 8'b00000000) && ((CC_COMPARADORCRASH_ALBERT_FROG_ROW_2_In_Bus | CC_COMPARADORCRASH_BACKGROUND_ROW_2_IN_BUS) == CC_COMPARADORCRASH_BACKGROUND_ROW_2_IN_BUS))
		CC_COMPARADORCRASH_Out_Bus = 2'b01;
	else if ((CC_COMPARADORCRASH_ALBERT_FROG_ROW_3_In_Bus != 8'b00000000) && ((CC_COMPARADORCRASH_ALBERT_FROG_ROW_3_In_Bus | CC_COMPARADORCRASH_BACKGROUND_ROW_3_IN_BUS) == CC_COMPARADORCRASH_BACKGROUND_ROW_3_IN_BUS))
		CC_COMPARADORCRASH_Out_Bus = 2'b01;
	else if ((CC_COMPARADORCRASH_ALBERT_FROG_ROW_4_In_Bus != 8'b00000000) && ((CC_COMPARADORCRASH_ALBERT_FROG_ROW_4_In_Bus | CC_COMPARADORCRASH_BACKGROUND_ROW_4_IN_BUS) == CC_COMPARADORCRASH_BACKGROUND_ROW_4_IN_BUS))
		CC_COMPARADORCRASH_Out_Bus = 2'b01;
	else if ((CC_COMPARADORCRASH_ALBERT_FROG_ROW_5_In_Bus != 8'b00000000) && ((CC_COMPARADORCRASH_ALBERT_FROG_ROW_5_In_Bus | CC_COMPARADORCRASH_BACKGROUND_ROW_5_IN_BUS) == CC_COMPARADORCRASH_BACKGROUND_ROW_5_IN_BUS))
		CC_COMPARADORCRASH_Out_Bus = 2'b01;
	else if ((CC_COMPARADORCRASH_ALBERT_FROG_ROW_6_In_Bus != 8'b00000000) && ((CC_COMPARADORCRASH_ALBERT_FROG_ROW_6_In_Bus | CC_COMPARADORCRASH_BACKGROUND_ROW_6_IN_BUS) == CC_COMPARADORCRASH_BACKGROUND_ROW_6_IN_BUS))
		CC_COMPARADORCRASH_Out_Bus = 2'b01;
	else if ((CC_COMPARADORCRASH_ALBERT_FROG_ROW_9_In_Bus != 8'b00000000) && ((CC_COMPARADORCRASH_ALBERT_FROG_ROW_9_In_Bus | CC_COMPARADORCRASH_BACKGROUND_ROW_9_IN_BUS) == CC_COMPARADORCRASH_BACKGROUND_ROW_9_IN_BUS))
		CC_COMPARADORCRASH_Out_Bus = 2'b01;
	else if ((CC_COMPARADORCRASH_ALBERT_FROG_ROW_10_In_Bus != 8'b00000000) && ((CC_COMPARADORCRASH_ALBERT_FROG_ROW_10_In_Bus | CC_COMPARADORCRASH_BACKGROUND_ROW_10_IN_BUS) == CC_COMPARADORCRASH_BACKGROUND_ROW_10_IN_BUS))
		CC_COMPARADORCRASH_Out_Bus = 2'b01;
	else if ((CC_COMPARADORCRASH_ALBERT_FROG_ROW_11_In_Bus != 8'b00000000) && ((CC_COMPARADORCRASH_ALBERT_FROG_ROW_11_In_Bus | CC_COMPARADORCRASH_BACKGROUND_ROW_11_IN_BUS) == CC_COMPARADORCRASH_BACKGROUND_ROW_11_IN_BUS))
		CC_COMPARADORCRASH_Out_Bus = 2'b01;	
	else if ((CC_COMPARADORCRASH_ALBERT_FROG_ROW_12_In_Bus != 8'b00000000) && ((CC_COMPARADORCRASH_ALBERT_FROG_ROW_12_In_Bus | CC_COMPARADORCRASH_BACKGROUND_ROW_12_IN_BUS) == CC_COMPARADORCRASH_BACKGROUND_ROW_12_IN_BUS))
		CC_COMPARADORCRASH_Out_Bus = 2'b01;
	else if ((CC_COMPARADORCRASH_ALBERT_FROG_ROW_13_In_Bus != 8'b00000000) && ((CC_COMPARADORCRASH_ALBERT_FROG_ROW_13_In_Bus | CC_COMPARADORCRASH_BACKGROUND_ROW_13_IN_BUS) == CC_COMPARADORCRASH_BACKGROUND_ROW_13_IN_BUS))
		CC_COMPARADORCRASH_Out_Bus = 2'b01;
	else if ((CC_COMPARADORCRASH_ALBERT_FROG_ROW_14_In_Bus != 8'b00000000) && ((CC_COMPARADORCRASH_ALBERT_FROG_ROW_14_In_Bus | CC_COMPARADORCRASH_END_GOAL_ROW_14_IN_BUS) == CC_COMPARADORCRASH_END_GOAL_ROW_14_IN_BUS))
		CC_COMPARADORCRASH_Out_Bus = 2'b01;
	else if ((CC_COMPARADORCRASH_ALBERT_FROG_ROW_14_In_Bus != 8'b00000000) && ((CC_COMPARADORCRASH_ALBERT_FROG_ROW_14_In_Bus | CC_COMPARADORCRASH_END_GOAL_ROW_14_IN_BUS) != CC_COMPARADORCRASH_END_GOAL_ROW_14_IN_BUS))
		CC_COMPARADORCRASH_Out_Bus = 2'b10;
	else 
		CC_COMPARADORCRASH_Out_Bus = 2'b00;
		
	if (CC_COMPARADORCRASH_ALBERT_FROG_ROW_7_In_Bus != 8'b00000000)
		CC_COMPARATORLOCATION_Out = 1'b1;
	else if (CC_COMPARADORCRASH_ALBERT_FROG_ROW_8_In_Bus != 8'b00000000)
		CC_COMPARATORLOCATION_Out = 1'b1;
	else if (CC_COMPARADORCRASH_ALBERT_FROG_ROW_9_In_Bus != 8'b00000000)
		CC_COMPARATORLOCATION_Out = 1'b1;
	else if (CC_COMPARADORCRASH_ALBERT_FROG_ROW_10_In_Bus != 8'b00000000)
		CC_COMPARATORLOCATION_Out = 1'b1;
	else if (CC_COMPARADORCRASH_ALBERT_FROG_ROW_11_In_Bus != 8'b00000000)
		CC_COMPARATORLOCATION_Out = 1'b1;
	else if (CC_COMPARADORCRASH_ALBERT_FROG_ROW_12_In_Bus != 8'b00000000)
		CC_COMPARATORLOCATION_Out = 1'b1;
	else if (CC_COMPARADORCRASH_ALBERT_FROG_ROW_13_In_Bus != 8'b00000000)
		CC_COMPARATORLOCATION_Out = 1'b1;
	else if (CC_COMPARADORCRASH_ALBERT_FROG_ROW_14_In_Bus != 8'b00000000)
		CC_COMPARATORLOCATION_Out = 1'b1;
	else
		CC_COMPARATORLOCATION_Out = 1'b0;

end

endmodule